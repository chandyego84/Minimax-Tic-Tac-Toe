module board(clk, rst, clr, en_player, en_cpu, selectPlayer[8:0], selectCPU[8:0],
    pos1, pos2, pos3, pos4, pos5, pos6, pos7, pos8, pos9);

input clk, rst, clr;


